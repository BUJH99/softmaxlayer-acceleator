/******************************************************************
* 모듈: ln_lut_exp (High-Precision) - Vivado 호환 최종 수정 버전
* 설명: ln(2) * exp 값을 저장하는 32-entry LUT (ROM)
* 포맷: 16-bit Signed Q4.11  (범위 ±16, 분해능 1/2048)
******************************************************************/
module ln_lut_exp (
    input  wire [4:0] addr,           // 5-bit 주소 (E = exp + 15)
    output reg  signed [15:0] data    // 16-bit Q4.11 형식
);
    always @(*) begin
        case (addr)
            // ★★★ 수정: 음수 부호를 숫자 리터럴 밖으로 빼서 단항 연산자로 사용 ★★★
            5'd0:  data = -16'sd21293; // E=0,  exp=-15, ≈ -10.396973
            5'd1:  data = -16'sd19874; // E=1,  exp=-14, ≈ -9.704102
            5'd2:  data = -16'sd18454; // E=2,  exp=-13, ≈ -9.010742
            5'd3:  data = -16'sd17035; // E=3,  exp=-12, ≈ -8.317871
            5'd4:  data = -16'sd15615; // E=4,  exp=-11, ≈ -7.624512
            5'd5:  data = -16'sd14196; // E=5,  exp=-10, ≈ -6.931641
            5'd6:  data = -16'sd12776; // E=6,  exp=-9,  ≈ -6.238281
            5'd7:  data = -16'sd11357; // E=7,  exp=-8,  ≈ -5.545410
            5'd8:  data = -16'sd9937;  // E=8,  exp=-7,  ≈ -4.852051
            5'd9:  data = -16'sd8517;  // E=9,  exp=-6,  ≈ -4.158691
            5'd10: data = -16'sd7098;  // E=10, exp=-5,  ≈ -3.465820
            5'd11: data = -16'sd5678;  // E=11, exp=-4,  ≈ -2.772461
            5'd12: data = -16'sd4259;  // E=12, exp=-3,  ≈ -2.079590
            5'd13: data = -16'sd2839;  // E=13, exp=-2,  ≈ -1.386230
            5'd14: data = -16'sd1420;  // E=14, exp=-1,  ≈ -0.693359
            5'd15: data = 16'sd0;      // E=15, exp=0,   ≈  0.000000
            5'd16: data = 16'sd1420;   // E=16, exp=+1,  ≈  0.693359
            5'd17: data = 16'sd2839;   // E=17, exp=+2,  ≈  1.386230
            5'd18: data = 16'sd4259;   // E=18, exp=+3,  ≈  2.079590
            5'd19: data = 16'sd5678;   // E=19, exp=+4,  ≈  2.772461
            5'd20: data = 16'sd7098;   // E=20, exp=+5,  ≈  3.465820
            5'd21: data = 16'sd8517;   // E=21, exp=+6,  ≈  4.158691
            5'd22: data = 16'sd9937;   // E=22, exp=+7,  ≈  4.852051
            5'd23: data = 16'sd11357;  // E=23, exp=+8,  ≈  5.545410
            5'd24: data = 16'sd12776;  // E=24, exp=+9,  ≈  6.238281
            5'd25: data = 16'sd14196;  // E=25, exp=+10, ≈  6.931641
            5'd26: data = 16'sd15615;  // E=26, exp=+11, ≈  7.624512
            5'd27: data = 16'sd17035;  // E=27, exp=+12, ≈  8.317871
            5'd28: data = 16'sd18454;  // E=28, exp=+13, ≈  9.010742
            5'd29: data = 16'sd19874;  // E=29, exp=+14, ≈  9.704102
            5'd30: data = 16'sd21293;  // E=30, exp=+15, ≈ 10.396973
            5'd31: data = 16'sd22713;  // E=31, exp=+16, ≈ 11.090332
            default: data = 16'sd0;
        endcase
    end
endmodule
