/******************************************************************
* 모듈: ln_lut_mant (High-Accuracy, Q0.16)
* 기능: y[a] = round( 65536 * ln(1 + a/256) ), a=0..255
* 포맷: 16-bit Unsigned Q0.16  (정밀도 극대화)
*
* 사용 맥락:
*   - mant(10b) = 정규화된 1.mant 의 소수부 상위 10비트
*   - addr = mant[9:2] (상위 8비트), frac = mant[1:0] (하위 2비트)
*   - 보간: y = y0 + ((y1 - y0) * frac) >>> 2
*     -> 근사 ln(1 + (addr + frac/4)/256)
*
* 검증 앵커:
*   - addr=  0: 0
*   - addr=128: ~26573 (≈ ln(1.5)*65536)
*   - addr=255: ~45298 (≈ ln(511/256)*65536)
******************************************************************/
module ln_lut_mant (
    input  wire [7:0]  addr,   // 8-bit 주소 (가수 상위 8비트)
    output reg  [15:0] data    // 16-bit Q0.16 (unsigned)
);
    always @(*) begin
        case (addr)
            8'd0: data = 16'd0;
            8'd1: data = 16'd256;
            8'd2: data = 16'd510;
            8'd3: data = 16'd764;
            8'd4: data = 16'd1016;
            8'd5: data = 16'd1268;
            8'd6: data = 16'd1518;
            8'd7: data = 16'd1768;
            8'd8: data = 16'd2017;
            8'd9: data = 16'd2264;
            8'd10: data = 16'd2511;
            8'd11: data = 16'd2757;
            8'd12: data = 16'd3002;
            8'd13: data = 16'd3246;
            8'd14: data = 16'd3489;
            8'd15: data = 16'd3732;
            8'd16: data = 16'd3973;
            8'd17: data = 16'd4214;
            8'd18: data = 16'd4453;
            8'd19: data = 16'd4692;
            8'd20: data = 16'd4929;
            8'd21: data = 16'd5166;
            8'd22: data = 16'd5401;
            8'd23: data = 16'd5636;
            8'd24: data = 16'd5869;
            8'd25: data = 16'd6102;
            8'd26: data = 16'd6334;
            8'd27: data = 16'd6564;
            8'd28: data = 16'd6794;
            8'd29: data = 16'd7023;
            8'd30: data = 16'd7251;
            8'd31: data = 16'd7478;
            8'd32: data = 16'd7704;
            8'd33: data = 16'd7929;
            8'd34: data = 16'd8154;
            8'd35: data = 16'd8377;
            8'd36: data = 16'd8600;
            8'd37: data = 16'd8821;
            8'd38: data = 16'd9042;
            8'd39: data = 16'd9262;
            8'd40: data = 16'd9481;
            8'd41: data = 16'd9699;
            8'd42: data = 16'd9916;
            8'd43: data = 16'd10133;
            8'd44: data = 16'd10348;
            8'd45: data = 16'd10563;
            8'd46: data = 16'd10777;
            8'd47: data = 16'd10990;
            8'd48: data = 16'd11202;
            8'd49: data = 16'd11413;
            8'd50: data = 16'd11624;
            8'd51: data = 16'd11833;
            8'd52: data = 16'd12042;
            8'd53: data = 16'd12250;
            8'd54: data = 16'd12457;
            8'd55: data = 16'd12663;
            8'd56: data = 16'd12868;
            8'd57: data = 16'd13073;
            8'd58: data = 16'd13276;
            8'd59: data = 16'd13479;
            8'd60: data = 16'd13681;
            8'd61: data = 16'd13882;
            8'd62: data = 16'd14082;
            8'd63: data = 16'd14282;
            8'd64: data = 16'd14480;
            8'd65: data = 16'd14678;
            8'd66: data = 16'd14875;
            8'd67: data = 16'd15071;
            8'd68: data = 16'd15266;
            8'd69: data = 16'd15460;
            8'd70: data = 16'd15654;
            8'd71: data = 16'd15847;
            8'd72: data = 16'd16039;
            8'd73: data = 16'd16230;
            8'd74: data = 16'd16420;
            8'd75: data = 16'd16610;
            8'd76: data = 16'd16798;
            8'd77: data = 16'd16986;
            8'd78: data = 16'd17173;
            8'd79: data = 16'd17359;
            8'd80: data = 16'd17545;
            8'd81: data = 16'd17729;
            8'd82: data = 16'd17913;
            8'd83: data = 16'd18096;
            8'd84: data = 16'd18278;
            8'd85: data = 16'd18459;
            8'd86: data = 16'd18639;
            8'd87: data = 16'd18819;
            8'd88: data = 16'd18998;
            8'd89: data = 16'd19176;
            8'd90: data = 16'd19353;
            8'd91: data = 16'd19530;
            8'd92: data = 16'd19705;
            8'd93: data = 16'd19880;
            8'd94: data = 16'd20055;
            8'd95: data = 16'd20228;
            8'd96: data = 16'd20400;
            8'd97: data = 16'd20572;
            8'd98: data = 16'd20743;
            8'd99: data = 16'd20913;
            8'd100: data = 16'd21082;
            8'd101: data = 16'd21251;
            8'd102: data = 16'd21419;
            8'd103: data = 16'd21586;
            8'd104: data = 16'd21753;
            8'd105: data = 16'd21919;
            8'd106: data = 16'd22084;
            8'd107: data = 16'd22248;
            8'd108: data = 16'd22412;
            8'd109: data = 16'd22575;
            8'd110: data = 16'd22737;
            8'd111: data = 16'd22899;
            8'd112: data = 16'd23060;
            8'd113: data = 16'd23220;
            8'd114: data = 16'd23380;
            8'd115: data = 16'd23539;
            8'd116: data = 16'd23697;
            8'd117: data = 16'd23855;
            8'd118: data = 16'd24012;
            8'd119: data = 16'd24168;
            8'd120: data = 16'd24324;
            8'd121: data = 16'd24479;
            8'd122: data = 16'd24633;
            8'd123: data = 16'd24787;
            8'd124: data = 16'd24940;
            8'd125: data = 16'd25092;
            8'd126: data = 16'd25244;
            8'd127: data = 16'd25395;
            8'd128: data = 16'd25545;
            8'd129: data = 16'd25695;
            8'd130: data = 16'd25843;
            8'd131: data = 16'd25992;
            8'd132: data = 16'd26139;
            8'd133: data = 16'd26286;
            8'd134: data = 16'd26433;
            8'd135: data = 16'd26578;
            8'd136: data = 16'd26723;
            8'd137: data = 16'd26868;
            8'd138: data = 16'd27012;
            8'd139: data = 16'd27155;
            8'd140: data = 16'd27298;
            8'd141: data = 16'd27440;
            8'd142: data = 16'd27581;
            8'd143: data = 16'd27722;
            8'd144: data = 16'd27862;
            8'd145: data = 16'd28002;
            8'd146: data = 16'd28141;
            8'd147: data = 16'd28279;
            8'd148: data = 16'd28417;
            8'd149: data = 16'd28554;
            8'd150: data = 16'd28691;
            8'd151: data = 16'd28827;
            8'd152: data = 16'd28963;
            8'd153: data = 16'd29098;
            8'd154: data = 16'd29232;
            8'd155: data = 16'd29366;
            8'd156: data = 16'd29499;
            8'd157: data = 16'd29632;
            8'd158: data = 16'd29764;
            8'd159: data = 16'd29895;
            8'd160: data = 16'd30026;
            8'd161: data = 16'd30156;
            8'd162: data = 16'd30286;
            8'd163: data = 16'd30415;
            8'd164: data = 16'd30544;
            8'd165: data = 16'd30672;
            8'd166: data = 16'd30800;
            8'd167: data = 16'd30927;
            8'd168: data = 16'd31053;
            8'd169: data = 16'd31179;
            8'd170: data = 16'd31305;
            8'd171: data = 16'd31430;
            8'd172: data = 16'd31554;
            8'd173: data = 16'd31678;
            8'd174: data = 16'd31802;
            8'd175: data = 16'd31924;
            8'd176: data = 16'd32047;
            8'd177: data = 16'd32168;
            8'd178: data = 16'd32290;
            8'd179: data = 16'd32410;
            8'd180: data = 16'd32530;
            8'd181: data = 16'd32650;
            8'd182: data = 16'd32769;
            8'd183: data = 16'd32887;
            8'd184: data = 16'd33005;
            8'd185: data = 16'd33123;
            8'd186: data = 16'd33239;
            8'd187: data = 16'd33356;
            8'd188: data = 16'd33471;
            8'd189: data = 16'd33586;
            8'd190: data = 16'd33701;
            8'd191: data = 16'd33815;
            8'd192: data = 16'd33928;
            8'd193: data = 16'd34041;
            8'd194: data = 16'd34154;
            8'd195: data = 16'd34266;
            8'd196: data = 16'd34377;
            8'd197: data = 16'd34488;
            8'd198: data = 16'd34598;
            8'd199: data = 16'd34708;
            8'd200: data = 16'd34817;
            8'd201: data = 16'd34926;
            8'd202: data = 16'd35034;
            8'd203: data = 16'd35142;
            8'd204: data = 16'd35249;
            8'd205: data = 16'd35356;
            8'd206: data = 16'd35462;
            8'd207: data = 16'd35568;
            8'd208: data = 16'd35673;
            8'd209: data = 16'd35778;
            8'd210: data = 16'd35882;
            8'd211: data = 16'd35986;
            8'd212: data = 16'd36089;
            8'd213: data = 16'd36192;
            8'd214: data = 16'd36294;
            8'd215: data = 16'd36395;
            8'd216: data = 16'd36497;
            8'd217: data = 16'd36597;
            8'd218: data = 16'd36697;
            8'd219: data = 16'd36797;
            8'd220: data = 16'd36896;
            8'd221: data = 16'd36995;
            8'd222: data = 16'd37093;
            8'd223: data = 16'd37191;
            8'd224: data = 16'd37288;
            8'd225: data = 16'd37385;
            8'd226: data = 16'd37481;
            8'd227: data = 16'd37577;
            8'd228: data = 16'd37673;
            8'd229: data = 16'd37768;
            8'd230: data = 16'd37862;
            8'd231: data = 16'd37956;
            8'd232: data = 16'd38050;
            8'd233: data = 16'd38143;
            8'd234: data = 16'd38235;
            8'd235: data = 16'd38327;
            8'd236: data = 16'd38419;
            8'd237: data = 16'd38510;
            8'd238: data = 16'd38600;
            8'd239: data = 16'd38691;
            8'd240: data = 16'd38780;
            8'd241: data = 16'd38869;
            8'd242: data = 16'd38958;
            8'd243: data = 16'd39046;
            8'd244: data = 16'd39134;
            8'd245: data = 16'd39222;
            8'd246: data = 16'd39309;
            8'd247: data = 16'd39395;
            8'd248: data = 16'd39481;
            8'd249: data = 16'd39567;
            8'd250: data = 16'd39652;
            8'd251: data = 16'd39737;
            8'd252: data = 16'd39821;
            8'd253: data = 16'd39905;
            8'd254: data = 16'd39988;
            8'd255: data = 16'd40071;
            
            default: data = 16'd0;
        endcase
    end
endmodule
